`include "add64bit.v"
`include "add1bit.v"

`timescale 1ns/1ps 
module add_64test;
reg signed [63:0] a;
reg signed [63:0] b;
wire signed [63:0] result;
wire overflow;
add64bit new(a,b,result,overflow);
initial begin
    $dumpfile("test_add64.vcd");
    $dumpvars(0,add_64test);
    a=64'b0000000000000000000000000000000000000000000000000000000000000000;
    b=64'b0000000000000000000000000000000000000000000000000000000000000000;
end

initial begin 
    $monitor("a=",a, " b= ",b," result =",result," overflow=",overflow);
    #5
    //add without overflow both positive numbers
    a=64'b1000000000000000000000000000000000000000000000000000000000000000;
    b=64'b0111111111111111111111111111111111111111111111111111111111111111;
    #5
    //add without overflow both negative numbers
    a=64'b1111111111111111111111111111111111111111111111111111111111111111;//-1
    b=64'b1111111111111111111111111111111111111111111111111111111111111011;//-5
    #5
    //add without overflow with positive and negative numbers
    a=64'b0000000000000000000000000000000000000000000000000000000000000001;//1
    b=64'b1111111111111111111111111111111111111111111111111111111111111011;//-5
    #5 
    //add with overflow with both positive numbers
    a=64'b0111111111111111111111111111111111111111111111111111111111111111;
    b=64'b0111111111111111111111111111111111111111111111111111111111111111;
    #5
    // add with overflow with both negative numbers
    a=64'b1000000000000000000000000000000000000000000000000000000000000000;
    b=64'b1000000000000000000000000000000000000000000000000000000000000001;
end
endmodule