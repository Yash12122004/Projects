`timescale 1ns / 1ps

module and1bit(c,a,b);
    input a,b;
    output c;
    and a1(c,a,b);
endmodule