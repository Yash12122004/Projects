`include "alu.v"
`timescale 1ns/1ps 

module alu_64test;

reg [1:0] control;
reg signed [63:0] a;
reg signed [63:0] b;
wire signed [63:0] result;
wire overflow;

alu new(control,a,b,result,overflow);

initial 
    begin 
        $dumpfile("alu_64test.vcd");
        $dumpvars(0,alu_64test);
        control=0;//add without overflow both positive numbers
        a=64'b1000000000000000000000000000000000000000000000000000000000000000;
        b=64'b0111111111111111111111111111111111111111111111111111111111111111;
    end

initial
    begin 
        $monitor(" control= ",control," a=",a, " b= ",b," result =",result," overflow=",overflow);
        //Add
        #5
        control=0;//add without overflow both negative numbers
        a=64'b1111111111111111111111111111111111111111111111111111111111111111;//-1
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;//-5
        #5
        control=0;//add without overflow with positive and negative numbers
        a=64'b0000000000000000000000000000000000000000000000000000000000000001;//1
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;//-5
        #5 
        control=0;//add with overflow with both positive numbers
        a=64'b0111111111111111111111111111111111111111111111111111111111111111;
        b=64'b0111111111111111111111111111111111111111111111111111111111111111;
        #5
        control=0;// add with overflow with both negative numbers
        a=64'b1000000000000000000000000000000000000000000000000000000000000000;
        b=64'b1000000000000000000000000000000000000000000000000000000000000001;
        
        //Sub
        #5 
        control=1;//sub without overflow with both positive numbers
        a=64'b0000000000000000000000000000000000000000000000000000000000000101;
        b=64'b0000000000000000000000000000000000000000000000000000000000000001;
        #5
        control=1;//sub without overflow with both negative numbers
        a=64'b1111111111111111111111111111111111111111111111111111111111111111;
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;
        #5
        control=1;//sub with overflow with positive and negative numbers
        a=64'b0111111111111111111111111111111111111111111111111111111111111111;
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;
        //And
        #5
        control=2;// and without overflow with both positive numbers;
        a=64'b0000000000000000000000000000000000000000000000000000000000000001;
        b=64'b0000000000000000000000000000000000000000000000000000000000000101;
        #5
        control=2;// and without overflow with both negative numbers;
        a=64'b1000000000000000000000000000000000000000000000000000000000000000;
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;
        #5
        control=2;// and without overflow with positive and negative numbers;
        a=64'b0111111111111111111111111111111111111111111111111111111111111111;
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;
        //Xor
        #5
        control=3;// xor without overflow with both positive numbers;
        a=64'b0000000000000000000000000000000000000000000000000000000000000001;
        b=64'b0000000000000000000000000000000000000000000000000000000000000101;
        #5
        control=3;// xor without overflow with both negative numbers;
        a=64'b1000000000000000000000000000000000000000000000000000000000000000;
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;
        #5
        control=3;// xor without overflow with positive and negative numbers;
        a=64'b0111111111111111111111111111111111111111111111111111111111111111;
        b=64'b1111111111111111111111111111111111111111111111111111111111111011;
        
    end
endmodule